module json112

[if debug]
fn log<T>(msg T) {
	println(msg)
}
