module vlsio
