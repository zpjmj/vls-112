module json112
