module json112

//后续添加utf16编码支持
fn utf16str_to_unicodepoint(str string, pos int) ?Unicode {
	return Unicode{}
}
