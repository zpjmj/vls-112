module meta

pub const (
	version = '0.0.1'
	description = 'V language simple server by 112'
)