// module tree2


// //二叉树
// struct Tree2{
// 	root int
// 	left_index
// 	left_tree Tree2
// 	right_index
// 	right_tree Tree2
// }

// pub fn (t Tree2) search(val int){

// 	if 	val <= t.root{
// 		if left_index.len == 0{
// 			return 
// 		}
// 		return t.left_tree.search(val)
// 	}else{
// 		if right_index.len == 0{
// 			return
// 		}
// 		return t.left_tree.search(val)
// 	}

// }








// pub fn

// fn  0 2
// ws  2 3
// name 3 7
// (  7 8
// )  8 9
// {  9 10
// ws 10 11
// name 11 12
// ( 12 13
// ) 13 14
// } 14 15
// {}fn 0 15
// ()fn 11 14






// fn main(){ a()}

// fn 


