module ast

pub struct JsonObject {
}
