module vlsio
