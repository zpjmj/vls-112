module json112